`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.01.2022 17:50:18
// Design Name: 
// Module Name: Data_RAM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module CONV1D_2nd_RAM
    #(
        Bit_width = 16,
        RAM_Depth = 44
    )
    (
        // Input
        input CLK,
        input Enable,
        input [4:0] Depth,
        input [3:0] Width,

        // Output
        output reg signed [Bit_width - 1 : 0] data_out_0,
        output reg signed [Bit_width - 1 : 0] data_out_1,
        output reg signed [Bit_width - 1 : 0] data_out_2,
        output reg signed [Bit_width - 1 : 0] data_out_3
    );

    // RAM reg creation
    (* RAM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_0 [0 : RAM_Depth - 1];
    (* RAM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_1 [0 : RAM_Depth - 1];
    (* RAM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_2 [0 : RAM_Depth - 1];
    (* RAM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_3 [0 : RAM_Depth - 1];

    always @ (negedge CLK) begin
        if (Enable) begin
            data_out_0 <= RAM_0[Width << 4 + Depth];
            data_out_1 <= RAM_1[Width << 4 + Depth];
            data_out_2 <= RAM_2[Width << 4 + Depth];
            data_out_3 <= RAM_3[Width << 4 + Depth];
        end else begin
            data_out_0 <= 0;
            data_out_1 <= 0;
            data_out_2 <= 0;
            data_out_3 <= 0;
        end
    end

    // Initialise the RAM
    initial begin
        RAM_0[0] = -16'd19;
        RAM_1[0] = 16'd6;
        RAM_2[0] = 16'd13;
        RAM_3[0] = 16'd3;
        RAM_0[1] = 16'd48;
        RAM_1[1] = 16'd0;
        RAM_2[1] = 16'd6;
        RAM_3[1] = -16'd22;
        RAM_0[2] = 16'd8;
        RAM_1[2] = 16'd10;
        RAM_2[2] = 16'd46;
        RAM_3[2] = 16'd27;
        RAM_0[3] = 16'd13;
        RAM_1[3] = -16'd1;
        RAM_2[3] = -16'd8;
        RAM_3[3] = -16'd27;
        RAM_0[4] = 16'd2;
        RAM_1[4] = 16'd4;
        RAM_2[4] = 16'd4;
        RAM_3[4] = -16'd23;
        RAM_0[5] = 16'd10;
        RAM_1[5] = -16'd11;
        RAM_2[5] = -16'd12;
        RAM_3[5] = -16'd21;
        RAM_0[6] = -16'd6;
        RAM_1[6] = -16'd15;
        RAM_2[6] = -16'd17;
        RAM_3[6] = 16'd36;
        RAM_0[7] = 16'd2;
        RAM_1[7] = -16'd7;
        RAM_2[7] = -16'd5;
        RAM_3[7] = -16'd7;
        RAM_0[8] = -16'd48;
        RAM_1[8] = 16'd4;
        RAM_2[8] = -16'd4;
        RAM_3[8] = 16'd23;
        RAM_0[9] = 16'd34;
        RAM_1[9] = 16'd2;
        RAM_2[9] = -16'd10;
        RAM_3[9] = -16'd14;
        RAM_0[10] = 16'd5;
        RAM_1[10] = -16'd11;
        RAM_2[10] = 16'd1;
        RAM_3[10] = 16'd18;
        RAM_0[11] = 16'd14;
        RAM_1[11] = 16'd18;
        RAM_2[11] = -16'd10;
        RAM_3[11] = -16'd35;
        RAM_0[12] = 16'd20;
        RAM_1[12] = -16'd7;
        RAM_2[12] = -16'd7;
        RAM_3[12] = 16'd6;
        RAM_0[13] = 16'd20;
        RAM_1[13] = -16'd26;
        RAM_2[13] = 16'd13;
        RAM_3[13] = 16'd5;
        RAM_0[14] = 16'd9;
        RAM_1[14] = -16'd7;
        RAM_2[14] = -16'd22;
        RAM_3[14] = 16'd4;
        RAM_0[15] = 16'd38;
        RAM_1[15] = -16'd17;
        RAM_2[15] = -16'd40;
        RAM_3[15] = 16'd2;
        RAM_0[4] = -16'd19;
        RAM_1[4] = -16'd2;
        RAM_2[4] = -16'd10;
        RAM_3[4] = -16'd15;
        RAM_0[5] = 16'd48;
        RAM_1[5] = 16'd9;
        RAM_2[5] = 16'd16;
        RAM_3[5] = 16'd10;
        RAM_0[6] = 16'd8;
        RAM_1[6] = -16'd9;
        RAM_2[6] = -16'd27;
        RAM_3[6] = -16'd49;
        RAM_0[7] = 16'd13;
        RAM_1[7] = 16'd36;
        RAM_2[7] = 16'd4;
        RAM_3[7] = 16'd22;
        RAM_0[8] = 16'd2;
        RAM_1[8] = 16'd11;
        RAM_2[8] = 16'd10;
        RAM_3[8] = 16'd15;
        RAM_0[9] = 16'd10;
        RAM_1[9] = 16'd13;
        RAM_2[9] = 16'd2;
        RAM_3[9] = 16'd13;
        RAM_0[10] = -16'd6;
        RAM_1[10] = -16'd2;
        RAM_2[10] = 16'd23;
        RAM_3[10] = -16'd19;
        RAM_0[11] = 16'd2;
        RAM_1[11] = -16'd4;
        RAM_2[11] = -16'd6;
        RAM_3[11] = -16'd4;
        RAM_0[12] = -16'd48;
        RAM_1[12] = -16'd4;
        RAM_2[12] = -16'd15;
        RAM_3[12] = 16'd2;
        RAM_0[13] = 16'd34;
        RAM_1[13] = 16'd6;
        RAM_2[13] = 16'd17;
        RAM_3[13] = -16'd19;
        RAM_0[14] = 16'd5;
        RAM_1[14] = -16'd2;
        RAM_2[14] = 16'd0;
        RAM_3[14] = -16'd17;
        RAM_0[15] = 16'd14;
        RAM_1[15] = -16'd4;
        RAM_2[15] = -16'd25;
        RAM_3[15] = 16'd19;
        RAM_0[16] = 16'd20;
        RAM_1[16] = -16'd19;
        RAM_2[16] = -16'd14;
        RAM_3[16] = -16'd16;
        RAM_0[17] = 16'd20;
        RAM_1[17] = -16'd35;
        RAM_2[17] = -16'd15;
        RAM_3[17] = -16'd8;
        RAM_0[18] = 16'd9;
        RAM_1[18] = -16'd19;
        RAM_2[18] = -16'd7;
        RAM_3[18] = -16'd7;
        RAM_0[19] = 16'd38;
        RAM_1[19] = 16'd17;
        RAM_2[19] = 16'd23;
        RAM_3[19] = 16'd53;
        RAM_0[8] = -16'd19;
        RAM_1[8] = 16'd26;
        RAM_2[8] = 16'd16;
        RAM_3[8] = 16'd4;
        RAM_0[9] = 16'd48;
        RAM_1[9] = 16'd2;
        RAM_2[9] = 16'd41;
        RAM_3[9] = -16'd15;
        RAM_0[10] = 16'd8;
        RAM_1[10] = -16'd25;
        RAM_2[10] = 16'd15;
        RAM_3[10] = -16'd54;
        RAM_0[11] = 16'd13;
        RAM_1[11] = -16'd45;
        RAM_2[11] = 16'd2;
        RAM_3[11] = 16'd4;
        RAM_0[12] = 16'd2;
        RAM_1[12] = 16'd20;
        RAM_2[12] = 16'd30;
        RAM_3[12] = -16'd39;
        RAM_0[13] = 16'd10;
        RAM_1[13] = -16'd33;
        RAM_2[13] = -16'd20;
        RAM_3[13] = 16'd21;
        RAM_0[14] = -16'd6;
        RAM_1[14] = 16'd43;
        RAM_2[14] = 16'd13;
        RAM_3[14] = 16'd22;
        RAM_0[15] = 16'd2;
        RAM_1[15] = 16'd24;
        RAM_2[15] = 16'd6;
        RAM_3[15] = 16'd0;
        RAM_0[16] = -16'd48;
        RAM_1[16] = 16'd4;
        RAM_2[16] = -16'd1;
        RAM_3[16] = 16'd7;
        RAM_0[17] = 16'd34;
        RAM_1[17] = -16'd4;
        RAM_2[17] = 16'd11;
        RAM_3[17] = 16'd12;
        RAM_0[18] = 16'd5;
        RAM_1[18] = 16'd15;
        RAM_2[18] = -16'd3;
        RAM_3[18] = -16'd21;
        RAM_0[19] = 16'd14;
        RAM_1[19] = 16'd75;
        RAM_2[19] = 16'd24;
        RAM_3[19] = -16'd31;
        RAM_0[20] = 16'd20;
        RAM_1[20] = -16'd2;
        RAM_2[20] = -16'd5;
        RAM_3[20] = -16'd4;
        RAM_0[21] = 16'd20;
        RAM_1[21] = 16'd44;
        RAM_2[21] = -16'd6;
        RAM_3[21] = 16'd5;
        RAM_0[22] = 16'd9;
        RAM_1[22] = -16'd25;
        RAM_2[22] = -16'd11;
        RAM_3[22] = 16'd4;
        RAM_0[23] = 16'd38;
        RAM_1[23] = -16'd45;
        RAM_2[23] = 16'd13;
        RAM_3[23] = 16'd54;
        RAM_0[12] = -16'd19;
        RAM_1[12] = 16'd5;
        RAM_2[12] = -16'd1;
        RAM_3[12] = -16'd12;
        RAM_0[13] = 16'd48;
        RAM_1[13] = 16'd15;
        RAM_2[13] = 16'd8;
        RAM_3[13] = -16'd39;
        RAM_0[14] = 16'd8;
        RAM_1[14] = 16'd27;
        RAM_2[14] = 16'd6;
        RAM_3[14] = 16'd13;
        RAM_0[15] = 16'd13;
        RAM_1[15] = 16'd34;
        RAM_2[15] = 16'd9;
        RAM_3[15] = 16'd7;
        RAM_0[16] = 16'd2;
        RAM_1[16] = 16'd7;
        RAM_2[16] = 16'd12;
        RAM_3[16] = 16'd22;
        RAM_0[17] = 16'd10;
        RAM_1[17] = -16'd20;
        RAM_2[17] = -16'd10;
        RAM_3[17] = -16'd15;
        RAM_0[18] = -16'd6;
        RAM_1[18] = -16'd16;
        RAM_2[18] = -16'd17;
        RAM_3[18] = -16'd15;
        RAM_0[19] = 16'd2;
        RAM_1[19] = -16'd15;
        RAM_2[19] = -16'd12;
        RAM_3[19] = -16'd9;
        RAM_0[20] = -16'd48;
        RAM_1[20] = -16'd2;
        RAM_2[20] = -16'd21;
        RAM_3[20] = 16'd39;
        RAM_0[21] = 16'd34;
        RAM_1[21] = 16'd27;
        RAM_2[21] = 16'd31;
        RAM_3[21] = -16'd35;
        RAM_0[22] = 16'd5;
        RAM_1[22] = 16'd2;
        RAM_2[22] = 16'd8;
        RAM_3[22] = -16'd21;
        RAM_0[23] = 16'd14;
        RAM_1[23] = -16'd7;
        RAM_2[23] = -16'd46;
        RAM_3[23] = -16'd36;
        RAM_0[24] = 16'd20;
        RAM_1[24] = -16'd6;
        RAM_2[24] = 16'd2;
        RAM_3[24] = 16'd22;
        RAM_0[25] = 16'd20;
        RAM_1[25] = -16'd46;
        RAM_2[25] = -16'd6;
        RAM_3[25] = -16'd7;
        RAM_0[26] = 16'd9;
        RAM_1[26] = -16'd26;
        RAM_2[26] = -16'd16;
        RAM_3[26] = 16'd35;
        RAM_0[27] = 16'd38;
        RAM_1[27] = -16'd11;
        RAM_2[27] = -16'd2;
        RAM_3[27] = 16'd1;
        RAM_0[16] = -16'd19;
        RAM_1[16] = -16'd6;
        RAM_2[16] = -16'd13;
        RAM_3[16] = -16'd18;
        RAM_0[17] = 16'd48;
        RAM_1[17] = 16'd19;
        RAM_2[17] = 16'd11;
        RAM_3[17] = -16'd33;
        RAM_0[18] = 16'd8;
        RAM_1[18] = 16'd9;
        RAM_2[18] = 16'd14;
        RAM_3[18] = -16'd2;
        RAM_0[19] = 16'd13;
        RAM_1[19] = 16'd14;
        RAM_2[19] = 16'd11;
        RAM_3[19] = 16'd6;
        RAM_0[20] = 16'd2;
        RAM_1[20] = 16'd5;
        RAM_2[20] = -16'd18;
        RAM_3[20] = 16'd11;
        RAM_0[21] = 16'd10;
        RAM_1[21] = -16'd2;
        RAM_2[21] = 16'd5;
        RAM_3[21] = 16'd13;
        RAM_0[22] = -16'd6;
        RAM_1[22] = -16'd24;
        RAM_2[22] = 16'd8;
        RAM_3[22] = 16'd1;
        RAM_0[23] = 16'd2;
        RAM_1[23] = -16'd20;
        RAM_2[23] = -16'd15;
        RAM_3[23] = -16'd6;
        RAM_0[24] = -16'd48;
        RAM_1[24] = -16'd10;
        RAM_2[24] = -16'd27;
        RAM_3[24] = 16'd18;
        RAM_0[25] = 16'd34;
        RAM_1[25] = 16'd13;
        RAM_2[25] = 16'd27;
        RAM_3[25] = -16'd39;
        RAM_0[26] = 16'd5;
        RAM_1[26] = -16'd4;
        RAM_2[26] = -16'd3;
        RAM_3[26] = -16'd20;
        RAM_0[27] = 16'd14;
        RAM_1[27] = -16'd27;
        RAM_2[27] = -16'd60;
        RAM_3[27] = 16'd45;
        RAM_0[28] = 16'd20;
        RAM_1[28] = -16'd15;
        RAM_2[28] = -16'd12;
        RAM_3[28] = -16'd7;
        RAM_0[29] = 16'd20;
        RAM_1[29] = -16'd59;
        RAM_2[29] = -16'd14;
        RAM_3[29] = 16'd28;
        RAM_0[30] = 16'd9;
        RAM_1[30] = -16'd16;
        RAM_2[30] = 16'd5;
        RAM_3[30] = 16'd28;
        RAM_0[31] = 16'd38;
        RAM_1[31] = 16'd37;
        RAM_2[31] = -16'd26;
        RAM_3[31] = -16'd9;
        RAM_0[20] = -16'd19;
        RAM_1[20] = -16'd9;
        RAM_2[20] = -16'd2;
        RAM_3[20] = -16'd15;
        RAM_0[21] = 16'd48;
        RAM_1[21] = 16'd32;
        RAM_2[21] = 16'd20;
        RAM_3[21] = 16'd36;
        RAM_0[22] = 16'd8;
        RAM_1[22] = 16'd13;
        RAM_2[22] = 16'd0;
        RAM_3[22] = -16'd25;
        RAM_0[23] = 16'd13;
        RAM_1[23] = 16'd54;
        RAM_2[23] = 16'd12;
        RAM_3[23] = 16'd27;
        RAM_0[24] = 16'd2;
        RAM_1[24] = 16'd13;
        RAM_2[24] = 16'd12;
        RAM_3[24] = 16'd14;
        RAM_0[25] = 16'd10;
        RAM_1[25] = 16'd21;
        RAM_2[25] = 16'd12;
        RAM_3[25] = 16'd7;
        RAM_0[26] = -16'd6;
        RAM_1[26] = -16'd15;
        RAM_2[26] = -16'd5;
        RAM_3[26] = 16'd1;
        RAM_0[27] = 16'd2;
        RAM_1[27] = -16'd30;
        RAM_2[27] = -16'd11;
        RAM_3[27] = -16'd9;
        RAM_0[28] = -16'd48;
        RAM_1[28] = -16'd8;
        RAM_2[28] = -16'd2;
        RAM_3[28] = -16'd1;
        RAM_0[29] = 16'd34;
        RAM_1[29] = 16'd28;
        RAM_2[29] = 16'd20;
        RAM_3[29] = 16'd1;
        RAM_0[30] = 16'd5;
        RAM_1[30] = -16'd21;
        RAM_2[30] = -16'd11;
        RAM_3[30] = 16'd2;
        RAM_0[31] = 16'd14;
        RAM_1[31] = -16'd29;
        RAM_2[31] = 16'd6;
        RAM_3[31] = 16'd6;
        RAM_0[32] = 16'd20;
        RAM_1[32] = -16'd17;
        RAM_2[32] = -16'd18;
        RAM_3[32] = -16'd23;
        RAM_0[33] = 16'd20;
        RAM_1[33] = -16'd45;
        RAM_2[33] = 16'd2;
        RAM_3[33] = 16'd15;
        RAM_0[34] = 16'd9;
        RAM_1[34] = -16'd3;
        RAM_2[34] = -16'd14;
        RAM_3[34] = -16'd15;
        RAM_0[35] = 16'd38;
        RAM_1[35] = 16'd1;
        RAM_2[35] = 16'd20;
        RAM_3[35] = -16'd10;
        RAM_0[24] = -16'd19;
        RAM_1[24] = 16'd21;
        RAM_2[24] = 16'd4;
        RAM_3[24] = 16'd2;
        RAM_0[25] = 16'd48;
        RAM_1[25] = 16'd11;
        RAM_2[25] = 16'd13;
        RAM_3[25] = 16'd9;
        RAM_0[26] = 16'd8;
        RAM_1[26] = -16'd4;
        RAM_2[26] = -16'd27;
        RAM_3[26] = -16'd20;
        RAM_0[27] = 16'd13;
        RAM_1[27] = -16'd34;
        RAM_2[27] = -16'd9;
        RAM_3[27] = -16'd40;
        RAM_0[28] = 16'd2;
        RAM_1[28] = -16'd42;
        RAM_2[28] = 16'd12;
        RAM_3[28] = 16'd4;
        RAM_0[29] = 16'd10;
        RAM_1[29] = -16'd6;
        RAM_2[29] = -16'd3;
        RAM_3[29] = 16'd44;
        RAM_0[30] = -16'd6;
        RAM_1[30] = -16'd9;
        RAM_2[30] = -16'd20;
        RAM_3[30] = 16'd7;
        RAM_0[31] = 16'd2;
        RAM_1[31] = 16'd5;
        RAM_2[31] = 16'd5;
        RAM_3[31] = 16'd21;
        RAM_0[32] = -16'd48;
        RAM_1[32] = 16'd8;
        RAM_2[32] = -16'd3;
        RAM_3[32] = 16'd5;
        RAM_0[33] = 16'd34;
        RAM_1[33] = 16'd5;
        RAM_2[33] = 16'd0;
        RAM_3[33] = -16'd50;
        RAM_0[34] = 16'd5;
        RAM_1[34] = 16'd22;
        RAM_2[34] = 16'd17;
        RAM_3[34] = 16'd31;
        RAM_0[35] = 16'd14;
        RAM_1[35] = 16'd83;
        RAM_2[35] = 16'd50;
        RAM_3[35] = 16'd10;
        RAM_0[36] = 16'd20;
        RAM_1[36] = 16'd8;
        RAM_2[36] = -16'd28;
        RAM_3[36] = -16'd27;
        RAM_0[37] = 16'd20;
        RAM_1[37] = 16'd67;
        RAM_2[37] = -16'd8;
        RAM_3[37] = -16'd3;
        RAM_0[38] = 16'd9;
        RAM_1[38] = -16'd1;
        RAM_2[38] = 16'd16;
        RAM_3[38] = 16'd13;
        RAM_0[39] = 16'd38;
        RAM_1[39] = -16'd76;
        RAM_2[39] = -16'd32;
        RAM_3[39] = -16'd14;
        RAM_0[28] = -16'd19;
        RAM_1[28] = -16'd11;
        RAM_2[28] = 16'd0;
        RAM_3[28] = 16'd0;
        RAM_0[29] = 16'd48;
        RAM_1[29] = 16'd16;
        RAM_2[29] = 16'd5;
        RAM_3[29] = -16'd23;
        RAM_0[30] = 16'd8;
        RAM_1[30] = 16'd55;
        RAM_2[30] = 16'd16;
        RAM_3[30] = -16'd2;
        RAM_0[31] = 16'd13;
        RAM_1[31] = -16'd10;
        RAM_2[31] = 16'd12;
        RAM_3[31] = -16'd15;
        RAM_0[32] = 16'd2;
        RAM_1[32] = 16'd5;
        RAM_2[32] = -16'd17;
        RAM_3[32] = -16'd18;
        RAM_0[33] = 16'd10;
        RAM_1[33] = -16'd9;
        RAM_2[33] = 16'd6;
        RAM_3[33] = 16'd10;
        RAM_0[34] = -16'd6;
        RAM_1[34] = -16'd29;
        RAM_2[34] = -16'd24;
        RAM_3[34] = 16'd13;
        RAM_0[35] = 16'd2;
        RAM_1[35] = -16'd16;
        RAM_2[35] = -16'd6;
        RAM_3[35] = 16'd5;
        RAM_0[36] = -16'd48;
        RAM_1[36] = -16'd22;
        RAM_2[36] = -16'd7;
        RAM_3[36] = 16'd16;
        RAM_0[37] = 16'd34;
        RAM_1[37] = 16'd11;
        RAM_2[37] = 16'd5;
        RAM_3[37] = -16'd7;
        RAM_0[38] = 16'd5;
        RAM_1[38] = 16'd6;
        RAM_2[38] = 16'd19;
        RAM_3[38] = 16'd24;
        RAM_0[39] = 16'd14;
        RAM_1[39] = -16'd26;
        RAM_2[39] = -16'd33;
        RAM_3[39] = 16'd3;
        RAM_0[40] = 16'd20;
        RAM_1[40] = -16'd8;
        RAM_2[40] = -16'd18;
        RAM_3[40] = -16'd1;
        RAM_0[41] = 16'd20;
        RAM_1[41] = -16'd30;
        RAM_2[41] = -16'd7;
        RAM_3[41] = -16'd11;
        RAM_0[42] = 16'd9;
        RAM_1[42] = 16'd13;
        RAM_2[42] = -16'd7;
        RAM_3[42] = -16'd1;
        RAM_0[43] = 16'd38;
        RAM_1[43] = -16'd24;
        RAM_2[43] = 16'd2;
        RAM_3[43] = -16'd28;
    end

endmodule